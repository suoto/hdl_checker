
entity entity_a is
end entity;

entity entity_a is
end entity;

entity entity_b is
end entity;
