
use work.entity_a;

use work.entity_b;

entity entity_c is
end entity;

architecture entity_c of entity_c is
begin
end entity_c;

