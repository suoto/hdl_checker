package sample_package is
end sample_package;
package body sample_package is
end sample_package;

